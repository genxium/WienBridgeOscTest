** Wien Bridge Oscillator No PWL with Diode Built-in Potential Kick-off and Stabilization 

* RC TUNING
R2	4	6	10K
C2	6 	3	16NF
R1	3 	0	10K
C1	3 	0	16NF
* NON-INVERTING OPAMP
R10	0	2	10K
R11	2	5	18K
XOP	3 2	4	OPAMP1
* AMPLITUDE STABILIZATION
R12	5	4	5K
D1	5	4	D1N914
D2	4	5	D1N914
*
.model	D1N914	D(Is=0.1p Rs=16 CJO=2p Tt=12n Bv=100 Ibv=0.1p)
*
* OPAMP MACRO MODEL, SINGLE-POLE 
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1      1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DC GAIN (100K) AND POLE 1 (100HZ)
EGAIN	3 0	1 2	100K
RP1	3	4	1K
CP1	4	0	1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
.ENDS

* ANALYSIS
** Without a PWL signal, the oscillation still starts but at a much later time!
.TRAN 	0.05MS 80MS
.CONTROL
RUN
PLOT	V(2) V(4) 
.ENDC
.END
