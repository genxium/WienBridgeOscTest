* OPAMP BASIC MATH MODEL POSITIVE FEEDBACK TESTING 

VIN 2 0 DC 0

XOP 1 2	3	OPAMP1
R1 0 1 1K 
R2 1 3 1K 

.SUBCKT OPAMP1      1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DC GAIN (100K) AND POLE 1 (100HZ)
EGAIN	3 0	1 2	100K
RP1	3	4	1K
CP1	4	0	1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
.ENDS

* DC Analysis
** .DC <srcname> <vstart> <vend> <vinc>
** ...
** .END

.DC VIN 0.25 5.0 0.25
.CONTROL
RUN
PLOT	V(2) V(3)
.ENDC
.END
