OPWIEN.CIR - OPAMP WIEN-BRIDGE OSCILLATOR
*
* CURRENT PULSE TO START OSCILLATIONS
IS	0	3	PWL(0US 0MA   10US 0.1MA   40US 0.1MA   50US 0MA   10MS 0MA)
*
* RC TUNING
R2	3	6	10K
C2	6 	0	16NF
R1	3 	4	10K
C1	3 	4	16NF
* NON-INVERTING OPAMP
R10	0	2	10K
R11	2	5	18K
XOP	3 2	4	OPAMP1
* AMPLITUDE STABILIZATION
R12	5	4	5K
D1	5	4	D1N914
D2	4	5	D1N914
*
.model	D1N914	D(Is=0.1p Rs=16 CJO=2p Tt=12n Bv=100 Ibv=0.1p)
*
* OPAMP MACRO MODEL, SINGLE-POLE 
* connections:      non-inverting input
*                   |   inverting input
*                   |   |   output
*                   |   |   |
.SUBCKT OPAMP1      1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DC GAIN (100K) AND POLE 1 (100HZ)
EGAIN	3 0	1 2	100K
RP1	3	4	1K
CP1	4	0	1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
.ENDS

* ANALYSIS
** No oscillation at all.
.TRAN 	0.05MS 100MS
.CONTROL
RUN
PLOT	V(4)
.ENDC
.END
