* OPAMP BASIC MATH MODEL MIXED FEEDBACK WITH DIODE BUILTIN POTENTIALS 

XOP 1 2	3	OPAMP1
R1 3 2 1K 
R2 2 0 1K 

R3 1 3 1K

D1	3	2 DIODE2	
D2	2	3 DIODE2	

.PARAM diodett=12n
.model	DIODE2	D(Is=0.1p Rs=16 CJO=2p Tt=diodett Bv=100 Ibv=0.1p)

.SUBCKT OPAMP1      1   2   6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DC GAIN (100K) AND POLE 1 (100HZ)
EGAIN	3 0	1 2	100K
RP1	3	4	1K
CP1	4	0	1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
.ENDS

* ANALYSIS
** There's an attenuating oscillation of V(2) which vanishes at around 25ns when diodett=12ns, which is apparently earlier than that of the `negative_feedback_with_diode_builtin_potentials` case.
.TRAN 	0.15NS 50NS
.CONTROL
RUN
PLOT	V(2) V(3)
.ENDC
.END
